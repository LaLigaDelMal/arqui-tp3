`timescale 1ns / 1ps


module Top_CPU(

    );
endmodule
