`timescale 1ns / 1ps
//Test bench top

module test_debug;

// Inputs
reg clk;
reg reset;
reg rx;


// Instantiate the module under test
TOP_TOP dut(
    clk,
    reset,
    rx
);

initial begin
    clk=0;
end

// Clock generation
always begin
    #5 clk = ~clk;
end

reg [9:0] load = 10'b1011011000;
reg [7:0] inst1[3:0];

integer i;
integer j;

initial begin
    inst1[0] = 8'b00111100;
    inst1[1] = 8'b00001000;
    inst1[2] = 8'b11111111;
    inst1[3] = 8'b11111111;

    i = 0;
    j = 0;
end

initial begin
    $display("Test debug");
    // RUN:  01110010
    // STEP: 01110011
    // LOAD: 01110011
    
    rx = 1;
    $display("Reset in progress");
    // Reset
    reset = 1;
    #10;
    reset = 0;
    
    $display("Reset Done");

    $display("Load");
    // lOAD
    
    // 104166
        
    for (i = 0; i < 10; i = i + 1) begin
        rx = load[i];
        $display("RX: %b", load[i]);
        #160;
    end

    	
    // Separar en 4 partes de 8 bits
    for (i = 0; i < 4; i = i + 1) begin
        rx = 0;
        #160;
        for (j = 0; j < 8; j = j + 1) begin
            rx = inst1[i][j];
            #160;
        end
        rx = 1;
        #160;
    end

    rx = 1;
    
    $display("Finish load");
    
    #300;
    $finish;
    
end



endmodule