`timescale 1ns / 1ps


module ID_EX_Reg(

    );
endmodule
