`timescale 1ns / 1ps


module Multiplexer(

    );
endmodule
