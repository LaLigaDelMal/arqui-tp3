`timescale 1ns / 1ps


module Debug_Unit(

    );
endmodule
