`timescale 1ns / 1ps


module Registers(

    );
endmodule
