`timescale 1ns / 1ps


module EX_MA_Reg(

    );
endmodule
