`timescale 1ns / 1ps


module Hazard_Unit(

    );
endmodule
