`timescale 1ns / 1ps


module CPU_Top(

    );
endmodule
