`timescale 1ns / 1ps


module MA_WB_Reg(

    );
endmodule
