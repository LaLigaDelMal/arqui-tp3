`timescale 1ns / 1ps


module Reg_MA_WB(

    );
endmodule
