`timescale 1ns / 1ps


module Forwarding_Unit(

    );
endmodule
