`timescale 1ns / 1ps


module IF_ID_Reg(

    );
endmodule
