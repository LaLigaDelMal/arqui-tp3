`timescale 1ns / 1ps


module Control_Unit(

    );
endmodule
